C6 - DIC  RTL INVERTER EXAMPLE
***CIRCUIT DESCRIPTION
VCC 6,0 DC 5
VIN 1,0 PULSE 0,5 2NS 2NS 2NS 80NS
RB1 1,2 10K
RC1 6,3 1K
Q1 3,2,0 QND
RB2 3,4 10K
Q2 5,4,0 QND
RC2 6,5 1K
*** OUTPUT SPEC:
.NP
.OUT V3 3,0 PRINT DC PLOT DC TRAN
.OUT V5 5,0 PRINT DC
***MODELS
.MODEL QND NPN BF=50 RB=70 RC=40 CCS=2PF TF=.1NS TR=10.NS CJE=.9PF
+  CJC=1.5PF PC=.85 VA=50
**** ANALYSIS
.TRAN 10NS 200NS 2NS 200NS
.SENS V3 V5
.DC VIN 0 5 .5
.END
  