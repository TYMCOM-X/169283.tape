.LIC 1  DIFFERENTIAL PAIR
***CIRCUIT:
VIN 1,0 AC 1 SIN 0 0.1 5MEG
VCC 8 0 DC 12
VEE 9,0 DC -12
Q1 4,2,6 QNL
Q2 5,3,6 QNL
RS1 1,2 1K
RS2 3,0 1K
RC1 4,8 10K
RC2 5,8 10K
Q3 6,7,9 QNL
Q4 7,7,9 QNL
RBIAS 7,8 20K
***OUTPUTS
.NP
.OUT V4 4,0 PRINT DC TRAN
.OUT V5 5,0 PRINT MAG PH DC TRAN PLOT MAG PH DC TRAN
***MODELS
.MODEL QNL NPN BF=80 RB=100 CCS=2PF TF=.3NS TR=6NS CJE=3PF CJC=2PF
+ VA=50
***ANALYSIS
.TRAN 10NS 500NS 1NS 500NS
.AC DEC 10 1 10GHZ
.DC VIN -.25 .25 .02
******
.END
 