.C5 - BRANCH CURRENT EXAMPLE
.NP 1
VS1 1,0 DC 10
VS2 3,0 DC 10
RS11 1,2 2
RS21 3,4 2
RS12 2,0 3
RS22 5,0 3
VCUR 4,5
.OUT ICAL VS1
.OUT ISHO VCUR
.DC 
.END
  