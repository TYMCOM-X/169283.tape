.C2 - SIMPLE RTL INVERTER
VCC 4,0 DC 5
VIN 1,0 PULSE 0,5,2NS 2NS 2NS 30NS
RB 1,2 10K
Q1 3,2,0 Q1
RC 4,3 1K
**** OUTPUT SPEC
.OUTPUT VC 3,0 PRINT DC PLOT TR 0 5
.NP
*** MODELS
.MODEL Q1 NPN BF=20 RB =100 TF=0.1NS CJC=2PF
*** ANALYSIS
.DC TC VIN 0,5 1
.TRAN 10NS 90NS 1NS 90NS
.END
