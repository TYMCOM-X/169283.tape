ONE TRANSIS AMP EXAMPLE
VCC 5 0 DC 12
VEE 6 0 DC -12
VIN 1 0 AC 1
RS 1 2 1K
Q1 3 2 4  X33
RC 5 3 500
RE 4 6 1K
CBY 4 0 1UFD
.OUT V3 3 0 PRINT MA PH
.DC OP
.SENSE V3
.AC DEC 10 1HZ TO 10MEGHZ
.MODEL X33 NPN BF=30 RB=50 VA=20
.END
 