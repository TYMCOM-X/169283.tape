. C1- SIMPLE DIFFERENTIAL PAIR
*** CIRCUIT DESCRIPTION:
VCC 7 0 DC 12
VEE 8,0 DC -12
VIN 1,0
RS1 1,2 1K
RS2 6,0 1K
Q1 3,2,4 MOD1
Q2 5,6,4 MOD1
RC1 7,3 10K
RC2 7,5 10K
RE 4,8 10K
*** DESCRIBE MODELS USED:
.MODEL MOD1 NPN BR=50 VA=50 IS=1.0E-12 RB=100
*** SPECIFY WHAT WE WISH TO OUTPUT:
.NP
.OUT VOUT 5,0  PLOT DC
*** WHAT TYPE OF ANALYSIS:
.DC TC VIN -1 5 .5
.END
 